** Profile: "SCHEMATIC1-simu_agua"  [ c:\users\joshu\onedrive\escritorio\modcomt\modulocomunicacion\simulaicionesorcad\simulacion_agua\simulacion_sensor_agua-pspicefiles\schematic1\simu_agua.sim ] 

** Creating circuit file "simu_agua.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/Cadence/SPB_17.4/tools/pspice/library/SS8050.lib" 
* From [PSPICE NETLIST] section of C:\Users\joshu\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 1000 1 10Meg
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
